module MIPS_TB();
wire		   	CLOCK_27;				//	27 MHz
reg		   	CLOCK_50=0;				//	50 MHz
wire			   EXT_CLOCK;				//	External Clock
////////////////////////	Push Button		////////////////////////
wire	   [3:0]	KEY;					//	Pushbutton[3:0]
////////////////////////	DPDT Switch		////////////////////////
reg	  [17:0]	SW;						//	Toggle Switch[17:0]
////////////////////////	7-SEG Dispaly	////////////////////////
wire	[6:0]	HEX0;					//	Seven Segment Digit 0
wire	[6:0]	HEX1;					//	Seven Segment Digit 1
wire	[6:0]	HEX2;					//	Seven Segment Digit 2
wire	[6:0]	HEX3;					//	Seven Segment Digit 3
wire	[6:0]	HEX4;					//	Seven Segment Digit 4
wire	[6:0]	HEX5;					//	Seven Segment Digit 5
wire	[6:0]	HEX6;					//	Seven Segment Digit 6
wire	[6:0]	HEX7;					//	Seven Segment Digit 7
////////////////////////////	LED		////////////////////////////
wire	[8:0]	LEDG;					//	LED Green[8:0]
wire  [17:0]	LEDR;					//	LED Red[17:0]
////////////////////////////	UART	////////////////////////////
//wire			UART_TXD;				//	UART Transmitter
//wire			   UART_RXD;				//	UART Receiver
////////////////////////////	IRDA	////////////////////////////
//wire			IRDA_TXD;				//	IRDA Transmitter
//wire			   IRDA_RXD;				//	IRDA Receiver
///////////////////////		SDRAM Interface	////////////////////////
wire	  [15:0]	DRAM_DQ;				//	SDRAM Data bus 16 Bits
wire  [11:0]	DRAM_ADDR;				//	SDRAM Address bus 12 Bits
wire			DRAM_LDQM;				//	SDRAM Low-byte Data Mask 
wire			DRAM_UDQM;				//	SDRAM High-byte Data Mask
wire			DRAM_WE_N;				//	SDRAM Write Enable
wire			DRAM_CAS_N;				//	SDRAM Column Address Strobe
wire			DRAM_RAS_N;				//	SDRAM Row Address Strobe
wire			DRAM_CS_N;				//	SDRAM Chip Select
wire			DRAM_BA_0;				//	SDRAM Bank Address 0
wire			DRAM_BA_1;				//	SDRAM Bank Address 0
wire			DRAM_CLK;				//	SDRAM Clock
wire			DRAM_CKE;				//	SDRAM Clock Enable
////////////////////////	Flash Interface	////////////////////////
wire	  [7:0]	FL_DQ;					//	FLASH Data bus 8 Bits
wire [21:0]	FL_ADDR;				//	FLASH Address bus 22 Bits
wire			FL_WE_N;				//	FLASH Write Enable
wire			FL_RST_N;				//	FLASH Reset
wire			FL_OE_N;				//	FLASH wire Enable
wire			FL_CE_N;				//	FLASH Chip Enable
////////////////////////	SRAM Interface	////////////////////////
wire	 [15:0]	SRAM_DQ;				//	SRAM Data bus 16 Bits
wire [17:0]	SRAM_ADDR;				//	SRAM Address bus 18 Bits
wire			SRAM_UB_N;				//	SRAM High-byte Data Mask 
wire			SRAM_LB_N;				//	SRAM Low-byte Data Mask 
wire			SRAM_WE_N;				//	SRAM Write Enable
wire			SRAM_CE_N;				//	SRAM Chip Enable
wire			SRAM_OE_N;				//	SRAM wire Enable
////////////////////	ISP1362 Interface	////////////////////////
wire	 [15:0]	OTG_DATA;				//	ISP1362 Data bus 16 Bits
wire  [1:0]	OTG_ADDR;				//	ISP1362 Address 2 Bits
wire			OTG_CS_N;				//	ISP1362 Chip Select
wire			OTG_RD_N;				//	ISP1362 Write
wire			OTG_WR_N;				//	ISP1362 Read
wire			OTG_RST_N;				//	ISP1362 Reset
wire			OTG_FSPEED;				//	USB Full Speed,	0 = Enable, Z = Disable
wire			OTG_LSPEED;				//	USB Low Speed, 	0 = Enable, Z = Disable
wire			   OTG_INT0;				//	ISP1362 Interrupt 0
wire			   OTG_INT1;				//	ISP1362 Interrupt 1
wire			   OTG_DREQ0;				//	ISP1362 DMA Request 0
wire			   OTG_DREQ1;				//	ISP1362 DMA Request 1
wire			OTG_DACK0_N;			//	ISP1362 DMA Acknowledge 0
wire			OTG_DACK1_N;			//	ISP1362 DMA Acknowledge 1
////////////////////	LCD Module 16X2	////////////////////////////
wire	  [7:0]	LCD_DATA;				//	LCD Data bus 8 bits
wire			LCD_ON;					//	LCD Power ON/OFF
wire			LCD_BLON;				//	LCD Back Light ON/OFF
wire			LCD_RW;					//	LCD Read/Write Select, 0 = Write, 1 = Read
wire			LCD_EN;					//	LCD Enable
wire			LCD_RS;					//	LCD Command/Data Select, 0 = Command, 1 = Data
////////////////////	SD Card Interface	////////////////////////
//wire	 [3:0]	SD_DAT;					//	SD Card Data
//wire			   SD_WP_N;				   //	SD write protect
//wire			   SD_CMD;					//	SD Card Command Signal
//wire			SD_CLK;					//	SD Card Clock
////////////////////////	I2C		////////////////////////////////
wire			   I2C_SDAT;				//	I2C Data
wire			I2C_SCLK;				//	I2C Clock
////////////////////////	PS2		////////////////////////////////
wire		 	   PS2_DAT;				//	PS2 Data
wire			   PS2_CLK;				//	PS2 Clock
////////////////////	USB JTAG link	////////////////////////////
wire  			TDI;					// CPLD -> FPGA (data in)
wire  			TCK;					// CPLD -> FPGA (clk)
wire  			TCS;					// CPLD -> FPGA (CS)
wire 			TDO;					// FPGA -> CPLD (data out)
////////////////////////	VGA			////////////////////////////
wire			VGA_CLK;   				//	VGA Clock
wire			VGA_HS;					//	VGA H_SYNC
wire			VGA_VS;					//	VGA V_SYNC
wire			VGA_BLANK;				//	VGA BLANK
wire			VGA_SYNC;				//	VGA SYNC
wire	[9:0]	VGA_R;   				//	VGA Red[9:0]
wire	[9:0]	VGA_G;	 				//	VGA Green[9:0]
wire	[9:0]	VGA_B;   				//	VGA Blue[9:0]
////////////////	Ethernet Interface	////////////////////////////
wire	[15:0]	ENET_DATA;				//	DM9000A DATA bus 16Bits
wire			ENET_CMD;				//	DM9000A Command/Data Select, 0 = Command, 1 = Data
wire			ENET_CS_N;				//	DM9000A Chip Select
wire			ENET_WR_N;				//	DM9000A Write
wire			ENET_RD_N;				//	DM9000A Read
wire			ENET_RST_N;				//	DM9000A Reset
wire			   ENET_INT;				//	DM9000A Interrupt
wire			ENET_CLK;				//	DM9000A Clock 25 MHz
////////////////////	Audio CODEC		////////////////////////////
wire			   AUD_ADCLRCK;			//	Audio CODEC ADC LR Clock
wire			   AUD_ADCDAT;				//	Audio CODEC ADC Data
wire			   AUD_DACLRCK;			//	Audio CODEC DAC LR Clock
wire			AUD_DACDAT;				//	Audio CODEC DAC Data
wire			   AUD_BCLK;				//	Audio CODEC Bit-Stream Clock
wire			AUD_XCK;				//	Audio CODEC Chip Clock
////////////////////	TV Devoder		////////////////////////////
wire	 [7:0]	TD_DATA;    			//	TV Decoder Data bus 8 bits
wire			   TD_HS;					//	TV Decoder H_SYNC
wire			   TD_VS;					//	TV Decoder V_SYNC
wire			TD_RESET;				//	TV Decoder Reset
wire          TD_CLK27;            //	TV Decoder 27MHz CLK
////////////////////////	GPIO	////////////////////////////////
wire	[35:0]	GPIO_0;					//	GPIO Connection 0
wire	[35:0]	GPIO_1;	
MIPS mips(
		////////////////////	Clock Input	 	////////////////////	 
		CLOCK_27,						//	27 MHz
		CLOCK_50,						//	50 MHz
		EXT_CLOCK,						//	External Clock
		////////////////////	Push Button		////////////////////
		KEY,							//	Pushbutton[3:0]
		////////////////////	DPDT Switch		////////////////////
		SW,								//	Toggle Switch[17:0]
		////////////////////	7-SEG Dispaly	////////////////////
		HEX0,							//	Seven Segment Digit 0
		HEX1,							//	Seven Segment Digit 1
		HEX2,							//	Seven Segment Digit 2
		HEX3,							//	Seven Segment Digit 3
		HEX4,							//	Seven Segment Digit 4
		HEX5,							//	Seven Segment Digit 5
		HEX6,							//	Seven Segment Digit 6
		HEX7,							//	Seven Segment Digit 7
		////////////////////////	LED		////////////////////////
		LEDG,							//	LED Green[8:0]
		LEDR,							//	LED Red[17:0]
		////////////////////////	UART	////////////////////////
		//UART_TXD,						//	UART Transmitter
		//UART_RXD,						//	UART Receiver
		////////////////////////	IRDA	////////////////////////
		//IRDA_TXD,						//	IRDA Transmitter
		//IRDA_RXD,						//	IRDA Receiver
		/////////////////////	SDRAM Interface		////////////////
		DRAM_DQ,						//	SDRAM Data bus 16 Bits
		DRAM_ADDR,						//	SDRAM Address bus 12 Bits
		DRAM_LDQM,						//	SDRAM Low-byte Data Mask 
		DRAM_UDQM,						//	SDRAM High-byte Data Mask
		DRAM_WE_N,						//	SDRAM Write Enable
		DRAM_CAS_N,						//	SDRAM Column Address Strobe
		DRAM_RAS_N,						//	SDRAM Row Address Strobe
		DRAM_CS_N,						//	SDRAM Chip Select
		DRAM_BA_0,						//	SDRAM Bank Address 0
		DRAM_BA_1,						//	SDRAM Bank Address 0
		DRAM_CLK,						//	SDRAM Clock
		DRAM_CKE,						//	SDRAM Clock Enable
		////////////////////	Flash Interface		////////////////
		FL_DQ,							//	FLASH Data bus 8 Bits
		FL_ADDR,						//	FLASH Address bus 22 Bits
		FL_WE_N,						//	FLASH Write Enable
		FL_RST_N,						//	FLASH Reset
		FL_OE_N,						//	FLASH Output Enable
		FL_CE_N,						//	FLASH Chip Enable
		////////////////////	SRAM Interface		////////////////
		SRAM_DQ,						//	SRAM Data bus 16 Bits
		SRAM_ADDR,						//	SRAM Address bus 18 Bits
		SRAM_UB_N,						//	SRAM High-byte Data Mask 
		SRAM_LB_N,						//	SRAM Low-byte Data Mask 
		SRAM_WE_N,						//	SRAM Write Enable
		SRAM_CE_N,						//	SRAM Chip Enable
		SRAM_OE_N,						//	SRAM Output Enable
		////////////////////	ISP1362 Interface	////////////////
		OTG_DATA,						//	ISP1362 Data bus 16 Bits
		OTG_ADDR,						//	ISP1362 Address 2 Bits
		OTG_CS_N,						//	ISP1362 Chip Select
		OTG_RD_N,						//	ISP1362 Write
		OTG_WR_N,						//	ISP1362 Read
		OTG_RST_N,						//	ISP1362 Reset
		OTG_FSPEED,						//	USB Full Speed,	0 = Enable, Z = Disable
		OTG_LSPEED,						//	USB Low Speed, 	0 = Enable, Z = Disable
		OTG_INT0,						//	ISP1362 Interrupt 0
		OTG_INT1,						//	ISP1362 Interrupt 1
		OTG_DREQ0,						//	ISP1362 DMA Request 0
		OTG_DREQ1,						//	ISP1362 DMA Request 1
		OTG_DACK0_N,					//	ISP1362 DMA Acknowledge 0
		OTG_DACK1_N,					//	ISP1362 DMA Acknowledge 1
		////////////////////	LCD Module 16X2		////////////////
		LCD_ON,							//	LCD Power ON/OFF
		LCD_BLON,						//	LCD Back Light ON/OFF
		LCD_RW,							//	LCD Read/Write Select, 0 = Write, 1 = Read
		LCD_EN,							//	LCD Enable
		LCD_RS,							//	LCD Command/Data Select, 0 = Command, 1 = Data
		LCD_DATA,						//	LCD Data bus 8 bits
		////////////////////	SD_Card Interface	////////////////
		//SD_DAT,							//	SD Card Data
		//SD_WP_N,						   //	SD Write protect 
		//SD_CMD,							//	SD Card Command Signal
		//SD_CLK,							//	SD Card Clock
		////////////////////	USB JTAG link	////////////////////
		TDI,  							// CPLD -> FPGA (data in)
		TCK,  							// CPLD -> FPGA (clk)
		TCS,  							// CPLD -> FPGA (CS)
	   TDO,  							// FPGA -> CPLD (data out)
		////////////////////	I2C		////////////////////////////
		I2C_SDAT,						//	I2C Data
		I2C_SCLK,						//	I2C Clock
		////////////////////	PS2		////////////////////////////
		PS2_DAT,						//	PS2 Data
		PS2_CLK,						//	PS2 Clock
		////////////////////	VGA		////////////////////////////
		VGA_CLK,   						//	VGA Clock
		VGA_HS,							//	VGA H_SYNC
		VGA_VS,							//	VGA V_SYNC
		VGA_BLANK,						//	VGA BLANK
		VGA_SYNC,						//	VGA SYNC
		VGA_R,   						//	VGA Red[9:0]
		VGA_G,	 						//	VGA Green[9:0]
		VGA_B,  						//	VGA Blue[9:0]
		////////////	Ethernet Interface	////////////////////////
		ENET_DATA,						//	DM9000A DATA bus 16Bits
		ENET_CMD,						//	DM9000A Command/Data Select, 0 = Command, 1 = Data
		ENET_CS_N,						//	DM9000A Chip Select
		ENET_WR_N,						//	DM9000A Write
		ENET_RD_N,						//	DM9000A Read
		ENET_RST_N,						//	DM9000A Reset
		ENET_INT,						//	DM9000A Interrupt
		ENET_CLK,						//	DM9000A Clock 25 MHz
		////////////////	Audio CODEC		////////////////////////
		AUD_ADCLRCK,					//	Audio CODEC ADC LR Clock
		AUD_ADCDAT,						//	Audio CODEC ADC Data
		AUD_DACLRCK,					//	Audio CODEC DAC LR Clock
		AUD_DACDAT,						//	Audio CODEC DAC Data
		AUD_BCLK,						//	Audio CODEC Bit-Stream Clock
		AUD_XCK,						//	Audio CODEC Chip Clock
		////////////////	TV Decoder		////////////////////////
		TD_DATA,    					//	TV Decoder Data bus 8 bits
		TD_HS,							//	TV Decoder H_SYNC
		TD_VS,							//	TV Decoder V_SYNC
		TD_RESET,						//	TV Decoder Reset
		TD_CLK27,                  //	TV Decoder 27MHz CLK
		////////////////////	GPIO	////////////////////////////
		GPIO_0,							//	GPIO Connection 0
		GPIO_1							//	GPIO Connection 1
	);
	initial repeat(500) 
	begin 
		#50 
		CLOCK_50 = ~CLOCK_50;
	end
	initial begin
		SW[0] = 1;
		#40
		SW[0] = 0;
	end
endmodule

